
`ifndef PKG_H
`define PKG_H
package pkg;
  import pkg_definitions::*;
  `include "simple_item_t.sv";
  `include "test_base_t.sv";
  `include "test1_t.sv";
  `include "test2_t.sv";
  `include "component_base_t.sv";
  `include "run_param_t.sv";
  `include "driver_t.sv";
  `include "collector_t.sv";
  `include "testbench_t.sv";
endpackage

`endif   