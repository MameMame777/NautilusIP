class sample_item;
  rand bit d,reset;
endclass