`define reg_addr1 32'h0000_0004
`define reg_addr2 32'h0000_0008